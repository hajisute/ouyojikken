`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   16:16:12 11/27/2018
// Design Name:   operation
// Module Name:   C:/Users/FPGA/Desktop/fpga-filter-hardware/operation_test.v
// Project Name:  memory
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: operation
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module operation_test_v;
	parameter PERIOD = 20;
	// Inputs
	reg [809:0] data_bus;
	reg clk;
	reg rst;
	reg refresh;

	// Outputs
	reg [9:0] out;
	wire [9:0] out_wire;
	always@(posedge clk)begin
		out <= out_wire;
	end
	// Instantiate the Unit Under Test (UUT)
	operation uut (
		.data_bus(data_bus), 
		.clk(clk), 
		.rst(rst), 
		.refresh(refresh), 
		.out(out_wire)
	);
	
	// �N���b�N�̐���


	initial begin
		// Initialize Inputs
		data_bus = 810'b000000000100000000110000000111000000111100000111110000000111000000001100000111110000000001000000001100000000010000000011000000011100000011110000011111000000011100000000110000011111000000000100000000110000000001000000001100000001110000001111000001111100000001110000000011000001111100000000010000000011000000000100000000110000000111000000111100000111110000000111000000001100000111110011111111001111111100111111110011111111001111111100111111110000011111000000011100000000110000011111000000000100000000110000000001000000001100000001110000001111000001111100000001110000000011000001111100000000010000000011000000000100000000110000000111000000111100000111110000000111000000001100000111110000000001000000001100000000010000000011000000011100000011110000011111000000011100000000110000011111000000000100000000110011111111;
		//000000000100000000110000000111000000111100000111110000000111000000001100000111110000000001000000001100000000010000000011000000011100000011110000011111000000011100000000110000011111000000000100000000110000000001000000001100000001110000001111000001111100000001110000000011000001111100000000010000000011000000000100000000110000000111000000111100000111110000000111000000001100000111110000000001000000001100000000010000000011000000011100000011110000011111000000011100000000110000011111000000000100000000110000000001000000001100000001110000001111000001111100000001110000000011000001111100000000010000000011000000000100000000110000000111000000111100000111110000000111000000001100000111110000000001000000001100000000010000000011000000011100000011110000011111000000011100000000110000011111000000000100000000110011111111;
		//111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		clk = 0;
		rst = 0;
		refresh = 0;

		// Wait 100 ns for global reset to finish
		// Add stimulus here

	end
	integer count = 0;
	   	// �N���b�N�̐���
	initial begin
	  clk = 1;
	  #(PERIOD / 4)
	  forever begin
		 #(PERIOD / 2) clk = 0;
		 #(PERIOD / 2) clk = 1;count = count + 1;
		 
	  end
	end
	// ���Z�b�g�̐���
	initial begin
	  rst = 1;
	  #(PERIOD * 2) rst = 0;
	end
      
endmodule

