`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    07:36:33 11/14/2018 
// Design Name: 
// Module Name:    medianfilter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module medianfilter#(
		//�e��f�l��bit���itag�i2b�j+��f�l�i8b�j�j
		parameter DATA_WIDTH = 8,
		parameter COLUMN_NUM = 7

	)(
		input wire clk,
		input wire rst,
		input wire refresh,
		input wire [DATA_WIDTH-1:0] in0,
		input wire [DATA_WIDTH-1:0] in1,
		input wire [DATA_WIDTH-1:0] in2,
		input wire [DATA_WIDTH-1:0] in3,
		input wire [DATA_WIDTH-1:0] in4,
		input wire [DATA_WIDTH-1:0] in5,
		input wire [DATA_WIDTH-1:0] in6,
		output reg [DATA_WIDTH-1:0] out
	);
	
	reg [8-1:0]input_tmp[7-1:0];//���͂��ꎞ�ۑ����邽�߂̃��W�X�^
	reg [8-1:0]queue_of_medians[7-1:0];//���͂̒����l��FIFO�ŋL�����郌�W�X�^
	wire [8-1:0]queue_of_medians_wire[7-1:0];//�����̃��W�X�^�̓��͗p���C��
	wire [8-1:0]out_wire;

	//sort_column:in0-6 -> out0-6(sorted)
	//sort_column�ȉ��͖������ł��B�B�B
	sort_column #(
		.DATA_WIDTH(DATA_WIDTH),
		.CULUMN_NUM(COLUMN_NUM)	  
	)sort_input(
		.clk(clk),
		.rst(rst),
		.in0(input_tmp[0]),
		.in1(input_tmp[1]),
		.in2(input_tmp[2]),
		.in3(input_tmp[3]),
		.in4(input_tmp[4]),
		.in5(input_tmp[5]),
		.in6(input_tmp[6]),	
		.out0(),
		.out1(),
		.out2(),
		.out3(queue_of_medians_wire[0]),
		.out4(),
		.out5(),
		.out6()

	);
	
	sort_column #(
		.DATA_WIDTH(DATA_WIDTH),
		.CULUMN_NUM(COLUMN_NUM)	  
	)sort_queue_of_medians(
		.clk(clk),
		.rst(rst),
		.in0(queue_of_medians[0]),
		.in1(queue_of_medians[1]),
		.in2(queue_of_medians[2]),
		.in3(queue_of_medians[3]),
		.in4(queue_of_medians[4]),
		.in5(queue_of_medians[5]),
		.in6(queue_of_medians[6]),
		.out0(),
		.out1(),
		.out2(),
		.out3(out_wire),
		.out4(),
		.out5(),
		.out6()		

	);


	integer i;
	
	always @(posedge clk) begin 
		if(rst|refresh)begin
			out <=  8'b00000000;
			for(i = 0; i < 7;i = i + 1)begin
				queue_of_medians[i] <= 8'b00000010;
				input_tmp[i] <= 8'b0;
			end
		end else begin
			out <= out_wire;
			queue_of_medians[0] <= queue_of_medians_wire[0];
			queue_of_medians[1] <= queue_of_medians_wire[1];
			queue_of_medians[2] <= queue_of_medians_wire[2];
			queue_of_medians[3] <= queue_of_medians_wire[3];
			queue_of_medians[4] <= queue_of_medians_wire[4];
			queue_of_medians[5] <= queue_of_medians_wire[5];
			queue_of_medians[6] <= queue_of_medians_wire[6];
			input_tmp[0] <= in0;
			input_tmp[1] <= in1;
			input_tmp[2] <= in2;
			input_tmp[3] <= in3;
			input_tmp[4] <= in4;
			input_tmp[5] <= in5;
			input_tmp[6] <= in6;
		end
	end

	assign queue_of_medians_wire[1] = queue_of_medians[0];
	assign queue_of_medians_wire[2] = queue_of_medians[1];
	assign queue_of_medians_wire[3] = queue_of_medians[2];
	assign queue_of_medians_wire[4] = queue_of_medians[3];
	assign queue_of_medians_wire[5] = queue_of_medians[4];
	assign queue_of_medians_wire[6] = queue_of_medians[5];
	

endmodule
